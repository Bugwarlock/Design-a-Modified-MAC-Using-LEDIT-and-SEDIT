* SPICE netlist written by S-Edit Win32 6.00
* Written on Oct 20, 2019 at 14:13:35

* Waveform probing commands
.probe
.options probefilename="two_Bits_FAdder."
+ probesdbfile="C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder.sdb"
+ probetopmodule="4_Bits_FAdder"

* No Ports in cell: PageID_Tanner
* End of module with no ports: PageID_Tanner

.SUBCKT Pad_Bond SIGNAL Subs
C1 SIGNAL Subs 0.25pF
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo, K.Schaefer  Oct 20, 2019  14:09:21
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module Pad_Bond / page Page0 
.ENDS

.SUBCKT PadBidirHE_2.0u DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
MN_4_1 OEB OE Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_2 N29 DataOut Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_3 N20 OE N29 Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_4 N29 OEB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_5 Pad N29 Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MN_4_6 DataInB DataInUnBuf Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MN_4_7 DataIn DataInB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
XPad_Bond_1 Pad Subs Pad_Bond
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Oct 20, 2019  14:09:21
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module PadBidirHE_2.0u / page Page0 
MP_4_1 OEB OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_2 N20 DataOut Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_3 N29 OEB N20 Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_4 N20 OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_5 Pad N20 Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MP_4_6 DataInB DataInUnBuf Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_7 DataIn DataInB Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
R1 Pad DataInUnBuf 100 TC1=0.0 TC2=0.0
.ENDS

.SUBCKT PadBidirHE DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
XPadBidirHE_2.0u_1 DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
+ PadBidirHE_2.0u
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Oct 20, 2019  14:09:21
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module PadBidirHE / page Page0 
.ENDS

.SUBCKT PadOut DataOut Pad Gnd Subs Vdd
XPadBidirHE_1 N6 N5 N4 DataOut Vdd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo  Oct 20, 2019  14:09:21
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module PadOut / page Page0 
.ENDS

.SUBCKT PadInC DataIn DataInB DataInUnBuf Pad Gnd Subs Vdd
XPadBidirHE_1 DataIn DataInB DataInUnBuf Gnd Gnd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Input Pad
* Designed by: D.Gunawan, J.Luo  Oct 20, 2019  14:08:07
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module PadInC / page Page0 
.ENDS

.SUBCKT XOR2 A B Out Gnd Vdd
M1 N2 B Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M2 N2 A Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M6 Out B N3 Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M5 N3 A Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M9 Out N2 Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
* Page Size:  5x7
* S-Edit  2-Input XOR Gate (TIB)
* Designed by: J. Luo  Oct 20, 2019  14:02:33
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module XOR2 / page Page0 
M3 N2 B N6 Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M4 N6 A Vdd Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M7 N5 A Vdd Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M10B Out N2 N5 Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M8 N4 B Vdd Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M10 Out N2 N4 Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
.ENDS

.SUBCKT NAND2 A B Out Gnd Vdd
M3 Out B 1 Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M4 1 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  2-Input NAND Gate (TIB)
* Designed by: J. Luo  Oct 20, 2019  14:02:33
* Schematic generated by S-Edit
* from file C:\Users\Mamad\Desktop\CA1-files\CA1\S-Edit\two_Bits_FAdder / module NAND2 / page Page0 
M2 Out B Vdd Vdd PMOS W='28*l' L='2*l' AS='144*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M1 Out A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
.ENDS

.SUBCKT 2_Bits_FAdder A B Cin Cout S Gnd Vdd
XNAND2_1 Cin N3 N5 Gnd Vdd NAND2
XNAND2_2 B A N6 Gnd Vdd NAND2
XNAND2_3 N6 N5 Cout Gnd Vdd NAND2
XXOR2_1 A B N3 Gnd Vdd XOR2
XXOR2_2 N3 Cin S Gnd Vdd XOR2
.ENDS

* Main circuit: 4_Bits_FAdder
X2_Bits_FAdder_1 N6 N7 N8 N10 N9 Gnd Vdd 2_Bits_FAdder
X2_Bits_FAdder_2 N1 N2 N3 N8 N4 Gnd Vdd 2_Bits_FAdder
X2_Bits_FAdder_3 N11 N12 N13 N3 N14 Gnd Vdd 2_Bits_FAdder
X2_Bits_FAdder_4 N16 N17 N18 N13 N19 Gnd Vdd 2_Bits_FAdder
XPadInC_1 N18 N20 N15 Cin Gnd Subs Vdd PadInC
XPadInC_2 N17 N23 N22 B1 Gnd Subs Vdd PadInC
XPadInC_3 N16 N27 N26 A1 Gnd Subs Vdd PadInC
XPadInC_4 N12 N31 N30 B2 Gnd Subs Vdd PadInC
XPadInC_5 N11 N33 N28 A2 Gnd Subs Vdd PadInC
XPadInC_6 N2 N38 N37 B3 Gnd Subs Vdd PadInC
XPadInC_7 N1 N35 N34 A3 Gnd Subs Vdd PadInC
XPadInC_8 N6 N41 N40 A4 Gnd Subs Vdd PadInC
XPadInC_9 N7 N44 N43 B4 Gnd Subs Vdd PadInC
XPadOut_1 N19 S1 Gnd Subs Vdd PadOut
XPadOut_2 N14 S2 Gnd Subs Vdd PadOut
XPadOut_3 N4 S3 Gnd Subs Vdd PadOut
XPadOut_4 N9 S4 Gnd Subs Vdd PadOut
XPadOut_5 N10 Cout Gnd Subs Vdd PadOut
* End of main circuit: 4_Bits_FAdder
